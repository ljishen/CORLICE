module corlice(led, sw);
   output [0:0] led;
   input [2:0] sw;

endmodule